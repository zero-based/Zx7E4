LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE timing IS
  -- Used for testbenches
  CONSTANT TIME_SPAN : TIME := 20 ns;
END PACKAGE;