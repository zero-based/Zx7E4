LIBRARY ieee;
LIBRARY vunit_lib;
USE ieee.std_logic_1164.ALL;
CONTEXT vunit_lib.vunit_context;

ENTITY register_file_tb IS
    GENERIC (runner_cfg : STRING);
END register_file_tb;

ARCHITECTURE tb OF register_file_tb IS

    CONSTANT COUNT_BITS : NATURAL := 5;
    CONSTANT REG_SIZE : NATURAL := 32;

    SIGNAL clk : std_logic;
    SIGNAL write_enable : std_logic;
    SIGNAL write_num : std_logic_vector (COUNT_BITS - 1 DOWNTO 0);
    SIGNAL read_num_1 : std_logic_vector (COUNT_BITS - 1 DOWNTO 0);
    SIGNAL read_num_2 : std_logic_vector (COUNT_BITS - 1 DOWNTO 0);
    SIGNAL write_data : std_logic_vector (REG_SIZE - 1 DOWNTO 0);
    SIGNAL read_data_1 : std_logic_vector (REG_SIZE - 1 DOWNTO 0);
    SIGNAL read_data_2 : std_logic_vector (REG_SIZE - 1 DOWNTO 0);

    TYPE test_case IS RECORD
        write_enable : std_logic;
        write_num : std_logic_vector (COUNT_BITS - 1 DOWNTO 0);
        read_num_1 : std_logic_vector (COUNT_BITS - 1 DOWNTO 0);
        read_num_2 : std_logic_vector (COUNT_BITS - 1 DOWNTO 0);
        write_data : std_logic_vector (REG_SIZE - 1 DOWNTO 0);
        read_data_1 : std_logic_vector (REG_SIZE - 1 DOWNTO 0);
        read_data_2 : std_logic_vector (REG_SIZE - 1 DOWNTO 0);
    END RECORD;

    TYPE test_case_array IS ARRAY (NATURAL RANGE <>) OF test_case;
    CONSTANT time_span : TIME := 1 us;

    CONSTANT test_cases : test_case_array := (
    -- Initial case
    ('0', "-----", "00000", "00001", "--------------------------------", "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU", "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"),

    -- Write/Read the same register
    ('1', "00000", "00000", "00000", "10101010101010101010101010101010", "10101010101010101010101010101010", "10101010101010101010101010101010"),

    -- Write/Read all Registers
    ('1', "00000", "-----", "-----", "00000000000000000000000000000001", "--------------------------------", "--------------------------------"),
    ('1', "00001", "-----", "-----", "00000000000000000000000000000010", "--------------------------------", "--------------------------------"),
    ('0', "-----", "00000", "00001", "--------------------------------", "00000000000000000000000000000001", "00000000000000000000000000000010"),
    
    ('1', "00010", "-----", "-----", "00000000000000000000000000000100", "--------------------------------", "--------------------------------"),
    ('1', "00011", "-----", "-----", "00000000000000000000000000001000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "00010", "00011", "--------------------------------", "00000000000000000000000000000100", "00000000000000000000000000001000"),

    ('1', "00100", "-----", "-----", "00000000000000000000000000010000", "--------------------------------", "--------------------------------"),
    ('1', "00101", "-----", "-----", "00000000000000000000000000100000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "00100", "00101", "--------------------------------", "00000000000000000000000000010000", "00000000000000000000000000100000"),
    
    ('1', "00110", "-----", "-----", "00000000000000000000000001000000", "--------------------------------", "--------------------------------"),
    ('1', "00111", "-----", "-----", "00000000000000000000000010000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "00110", "00111", "--------------------------------", "00000000000000000000000001000000", "00000000000000000000000010000000"),
    
    ('1', "01000", "-----", "-----", "00000000000000000000000100000000", "--------------------------------", "--------------------------------"),
    ('1', "01001", "-----", "-----", "00000000000000000000001000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "01000", "01001", "--------------------------------", "00000000000000000000000100000000", "00000000000000000000001000000000"),
    
    ('1', "01010", "-----", "-----", "00000000000000000000010000000000", "--------------------------------", "--------------------------------"),
    ('1', "01011", "-----", "-----", "00000000000000000000100000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "01010", "01011", "--------------------------------", "00000000000000000000010000000000", "00000000000000000000100000000000"),

    ('1', "01100", "-----", "-----", "00000000000000000001000000000000", "--------------------------------", "--------------------------------"),
    ('1', "01101", "-----", "-----", "00000000000000000010000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "01100", "01101", "--------------------------------", "00000000000000000001000000000000", "00000000000000000010000000000000"),

    ('1', "01110", "-----", "-----", "00000000000000000100000000000000", "--------------------------------", "--------------------------------"),
    ('1', "01111", "-----", "-----", "00000000000000001000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "01110", "01111", "--------------------------------", "00000000000000000100000000000000", "00000000000000001000000000000000"),

    ('1', "10000", "-----", "-----", "00000000000000010000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "10001", "-----", "-----", "00000000000000100000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "10000", "10001", "--------------------------------", "00000000000000010000000000000000", "00000000000000100000000000000000"),

    ('1', "10010", "-----", "-----", "00000000000001000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "10011", "-----", "-----", "00000000000010000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "10010", "10011", "--------------------------------", "00000000000001000000000000000000", "00000000000010000000000000000000"),

    ('1', "10100", "-----", "-----", "00000000000100000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "10101", "-----", "-----", "00000000001000000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "10100", "10101", "--------------------------------", "00000000000100000000000000000000", "00000000001000000000000000000000"),

    ('1', "10110", "-----", "-----", "00000000010000000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "10111", "-----", "-----", "00000000100000000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "10110", "10111", "--------------------------------", "00000000010000000000000000000000", "00000000100000000000000000000000"),

    ('1', "11000", "-----", "-----", "00000001000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "11001", "-----", "-----", "00000010000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "11000", "11001", "--------------------------------", "00000001000000000000000000000000", "00000010000000000000000000000000"),

    ('1', "11010", "-----", "-----", "00000100000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "11011", "-----", "-----", "00001000000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "11010", "11011", "--------------------------------", "00000100000000000000000000000000", "00001000000000000000000000000000"),

    ('1', "11100", "-----", "-----", "00010000000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "11101", "-----", "-----", "00100000000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "11100", "11101", "--------------------------------", "00010000000000000000000000000000", "00100000000000000000000000000000"),
    
    ('1', "11110", "-----", "-----", "01000000000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('1', "11111", "-----", "-----", "10000000000000000000000000000000", "--------------------------------", "--------------------------------"),
    ('0', "-----", "11110", "11111", "--------------------------------", "01000000000000000000000000000000", "10000000000000000000000000000000")
    );

BEGIN

    UUT : ENTITY work.register_file GENERIC MAP (
        COUNT_BITS => COUNT_BITS,
        REG_SIZE => REG_SIZE
        )
        PORT MAP(
            clk => clk,
            write_enable => write_enable,
            write_num => write_num,
            read_num_1 => read_num_1,
            read_num_2 => read_num_2,
            write_data => write_data,
            read_data_1 => read_data_1,
            read_data_2 => read_data_2
        );

    clk_process : PROCESS
    BEGIN
        clk <= '0';
        WAIT FOR time_span/2;
        clk <= '1';
        WAIT FOR time_span/2;
    END PROCESS;

    main : PROCESS
    BEGIN
        test_runner_setup(runner, runner_cfg);

        FOR i IN test_cases'RANGE LOOP

            write_enable <= test_cases(i).write_enable;
            write_num <= test_cases(i).write_num;
            read_num_1 <= test_cases(i).read_num_1;
            read_num_2 <= test_cases(i).read_num_2;
            write_data <= test_cases(i).write_data;

            WAIT FOR time_span;
            ASSERT (read_data_1 = test_cases(i).read_data_1 or test_cases(i).read_data_1 = "--------------------------------")
            REPORT "test " & INTEGER'image(i) & " failed [Read Data 1]" SEVERITY error;
            ASSERT (read_data_2 = test_cases(i).read_data_2 or test_cases(i).read_data_2 = "--------------------------------")
            REPORT "test " & INTEGER'image(i) & " failed [Read Data 2]" SEVERITY error;

        END LOOP;

        WAIT FOR time_span;
        test_runner_cleanup(runner);
        WAIT;

    END PROCESS;

END tb;