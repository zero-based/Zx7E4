LIBRARY ieee;
LIBRARY vunit_lib;
USE ieee.std_logic_1164.ALL;
USE work.timing.ALL;
CONTEXT vunit_lib.vunit_context;

ENTITY register_file_tb IS
  GENERIC (runner_cfg : STRING);
END register_file_tb;

ARCHITECTURE tb OF register_file_tb IS

  CONSTANT N : NATURAL := 5;
  CONSTANT SIZE : NATURAL := 32;

  TYPE test_t IS RECORD
    wr_ena : std_logic;
    wr_sel : std_logic_vector (N - 1 DOWNTO 0);
    rd_sel_1 : std_logic_vector (N - 1 DOWNTO 0);
    rd_sel_2 : std_logic_vector (N - 1 DOWNTO 0);
    wr : std_logic_vector (SIZE - 1 DOWNTO 0);
    rd_1 : std_logic_vector (SIZE - 1 DOWNTO 0);
    rd_2 : std_logic_vector (SIZE - 1 DOWNTO 0);
  END RECORD;

  TYPE test_array_t IS ARRAY (NATURAL RANGE <>) OF test_t;

  SIGNAL clk : std_logic;
  SIGNAL sig : test_t;

  CONSTANT tests : test_array_t := (
  -- Initial case
  ('0', "-----", "00000", "00001", "--------------------------------", "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU", "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"),

  -- Write/Read the same register
  ('1', "00000", "00000", "00000", "10101010101010101010101010101010", "10101010101010101010101010101010", "10101010101010101010101010101010"),

  -- Write/Read all Registers
  ('1', "00000", "-----", "-----", "00000000000000000000000000000001", "--------------------------------", "--------------------------------"),
  ('1', "00001", "-----", "-----", "00000000000000000000000000000010", "--------------------------------", "--------------------------------"),
  ('0', "-----", "00000", "00001", "--------------------------------", "00000000000000000000000000000001", "00000000000000000000000000000010"),

  ('1', "00010", "-----", "-----", "00000000000000000000000000000100", "--------------------------------", "--------------------------------"),
  ('1', "00011", "-----", "-----", "00000000000000000000000000001000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "00010", "00011", "--------------------------------", "00000000000000000000000000000100", "00000000000000000000000000001000"),

  ('1', "00100", "-----", "-----", "00000000000000000000000000010000", "--------------------------------", "--------------------------------"),
  ('1', "00101", "-----", "-----", "00000000000000000000000000100000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "00100", "00101", "--------------------------------", "00000000000000000000000000010000", "00000000000000000000000000100000"),

  ('1', "00110", "-----", "-----", "00000000000000000000000001000000", "--------------------------------", "--------------------------------"),
  ('1', "00111", "-----", "-----", "00000000000000000000000010000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "00110", "00111", "--------------------------------", "00000000000000000000000001000000", "00000000000000000000000010000000"),

  ('1', "01000", "-----", "-----", "00000000000000000000000100000000", "--------------------------------", "--------------------------------"),
  ('1', "01001", "-----", "-----", "00000000000000000000001000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "01000", "01001", "--------------------------------", "00000000000000000000000100000000", "00000000000000000000001000000000"),

  ('1', "01010", "-----", "-----", "00000000000000000000010000000000", "--------------------------------", "--------------------------------"),
  ('1', "01011", "-----", "-----", "00000000000000000000100000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "01010", "01011", "--------------------------------", "00000000000000000000010000000000", "00000000000000000000100000000000"),

  ('1', "01100", "-----", "-----", "00000000000000000001000000000000", "--------------------------------", "--------------------------------"),
  ('1', "01101", "-----", "-----", "00000000000000000010000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "01100", "01101", "--------------------------------", "00000000000000000001000000000000", "00000000000000000010000000000000"),

  ('1', "01110", "-----", "-----", "00000000000000000100000000000000", "--------------------------------", "--------------------------------"),
  ('1', "01111", "-----", "-----", "00000000000000001000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "01110", "01111", "--------------------------------", "00000000000000000100000000000000", "00000000000000001000000000000000"),

  ('1', "10000", "-----", "-----", "00000000000000010000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "10001", "-----", "-----", "00000000000000100000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "10000", "10001", "--------------------------------", "00000000000000010000000000000000", "00000000000000100000000000000000"),

  ('1', "10010", "-----", "-----", "00000000000001000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "10011", "-----", "-----", "00000000000010000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "10010", "10011", "--------------------------------", "00000000000001000000000000000000", "00000000000010000000000000000000"),

  ('1', "10100", "-----", "-----", "00000000000100000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "10101", "-----", "-----", "00000000001000000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "10100", "10101", "--------------------------------", "00000000000100000000000000000000", "00000000001000000000000000000000"),

  ('1', "10110", "-----", "-----", "00000000010000000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "10111", "-----", "-----", "00000000100000000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "10110", "10111", "--------------------------------", "00000000010000000000000000000000", "00000000100000000000000000000000"),

  ('1', "11000", "-----", "-----", "00000001000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "11001", "-----", "-----", "00000010000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "11000", "11001", "--------------------------------", "00000001000000000000000000000000", "00000010000000000000000000000000"),

  ('1', "11010", "-----", "-----", "00000100000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "11011", "-----", "-----", "00001000000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "11010", "11011", "--------------------------------", "00000100000000000000000000000000", "00001000000000000000000000000000"),

  ('1', "11100", "-----", "-----", "00010000000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "11101", "-----", "-----", "00100000000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "11100", "11101", "--------------------------------", "00010000000000000000000000000000", "00100000000000000000000000000000"),

  ('1', "11110", "-----", "-----", "01000000000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('1', "11111", "-----", "-----", "10000000000000000000000000000000", "--------------------------------", "--------------------------------"),
  ('0', "-----", "11110", "11111", "--------------------------------", "01000000000000000000000000000000", "10000000000000000000000000000000")
  );

BEGIN

  UUT : ENTITY work.register_file GENERIC MAP (
    N => N,
    SIZE => SIZE
    )
    PORT MAP(
      clk => clk,
      wr_ena => sig.wr_ena,
      wr_sel => sig.wr_sel,
      rd_sel_1 => sig.rd_sel_1,
      rd_sel_2 => sig.rd_sel_2,
      wr => sig.wr,
      rd_1 => sig.rd_1,
      rd_2 => sig.rd_2
    );

  tick : PROCESS
  BEGIN
    clk <= '0';
    WAIT FOR TIME_SPAN / 2;
    clk <= '1';
    WAIT FOR TIME_SPAN / 2;
  END PROCESS;

  main : PROCESS
  BEGIN
    test_runner_setup(runner, runner_cfg);

    FOR i IN tests'RANGE LOOP

      sig.wr_ena <= tests(i).wr_ena;
      sig.wr_sel <= tests(i).wr_sel;
      sig.rd_sel_1 <= tests(i).rd_sel_1;
      sig.rd_sel_2 <= tests(i).rd_sel_2;
      sig.wr <= tests(i).wr;

      WAIT FOR TIME_SPAN;

      ASSERT (sig.rd_1 = tests(i).rd_1 OR tests(i).rd_1 = "--------------------------------")
      REPORT "test " & INTEGER'image(i) & " failed [rd_1]" SEVERITY error;

      ASSERT (sig.rd_2 = tests(i).rd_2 OR tests(i).rd_2 = "--------------------------------")
      REPORT "test " & INTEGER'image(i) & " failed [rd_2]" SEVERITY error;

    END LOOP;

    WAIT FOR TIME_SPAN;
    test_runner_cleanup(runner);
    WAIT;

  END PROCESS;

END tb;