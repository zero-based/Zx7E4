LIBRARY ieee;
LIBRARY vunit_lib;
USE ieee.std_logic_1164.ALL;
USE work.timing.ALL;
CONTEXT vunit_lib.vunit_context;

ENTITY register_file_tb IS
  GENERIC (runner_cfg : STRING);
END register_file_tb;

ARCHITECTURE tb OF register_file_tb IS

  CONSTANT N : NATURAL := 5;
  CONSTANT SIZE : NATURAL := 32;

  TYPE test_t IS RECORD
    wr_ena : std_logic;
    wr_sel : std_logic_vector (N - 1 DOWNTO 0);
    rd_sel_1 : std_logic_vector (N - 1 DOWNTO 0);
    rd_sel_2 : std_logic_vector (N - 1 DOWNTO 0);
    wr : std_logic_vector (SIZE - 1 DOWNTO 0);
    rd_1 : std_logic_vector (SIZE - 1 DOWNTO 0);
    rd_2 : std_logic_vector (SIZE - 1 DOWNTO 0);
  END RECORD;

  TYPE test_array_t IS ARRAY (NATURAL RANGE <>) OF test_t;

  SIGNAL clk : std_logic;
  SIGNAL sig : test_t;

  CONSTANT tests : test_array_t := (
  -- Initial case
  ('0', "-----", "00000", "00001", X"--------", X"UUUUUUUU", X"UUUUUUUU"),

  -- Write/Read the same register
  ('1', "00000", "00000", "00000", X"AAAAAAAA", X"AAAAAAAA", X"AAAAAAAA"),

  -- Write/Read all Registers
  ('1', "00000", "-----", "-----", X"00000001", X"--------", X"--------"),
  ('1', "00001", "-----", "-----", X"00000002", X"--------", X"--------"),
  ('0', "-----", "00000", "00001", X"--------", X"00000001", X"00000002"),

  ('1', "00010", "-----", "-----", X"00000004", X"--------", X"--------"),
  ('1', "00011", "-----", "-----", X"00000008", X"--------", X"--------"),
  ('0', "-----", "00010", "00011", X"--------", X"00000004", X"00000008"),

  ('1', "00100", "-----", "-----", X"00000010", X"--------", X"--------"),
  ('1', "00101", "-----", "-----", X"00000020", X"--------", X"--------"),
  ('0', "-----", "00100", "00101", X"--------", X"00000010", X"00000020"),

  ('1', "00110", "-----", "-----", X"00000040", X"--------", X"--------"),
  ('1', "00111", "-----", "-----", X"00000080", X"--------", X"--------"),
  ('0', "-----", "00110", "00111", X"--------", X"00000040", X"00000080"),

  ('1', "01000", "-----", "-----", X"00000100", X"--------", X"--------"),
  ('1', "01001", "-----", "-----", X"00000200", X"--------", X"--------"),
  ('0', "-----", "01000", "01001", X"--------", X"00000100", X"00000200"),

  ('1', "01010", "-----", "-----", X"00000400", X"--------", X"--------"),
  ('1', "01011", "-----", "-----", X"00000800", X"--------", X"--------"),
  ('0', "-----", "01010", "01011", X"--------", X"00000400", X"00000800"),

  ('1', "01100", "-----", "-----", X"00001000", X"--------", X"--------"),
  ('1', "01101", "-----", "-----", X"00002000", X"--------", X"--------"),
  ('0', "-----", "01100", "01101", X"--------", X"00001000", X"00002000"),

  ('1', "01110", "-----", "-----", X"00004000", X"--------", X"--------"),
  ('1', "01111", "-----", "-----", X"00008000", X"--------", X"--------"),
  ('0', "-----", "01110", "01111", X"--------", X"00004000", X"00008000"),

  ('1', "10000", "-----", "-----", X"00010000", X"--------", X"--------"),
  ('1', "10001", "-----", "-----", X"00020000", X"--------", X"--------"),
  ('0', "-----", "10000", "10001", X"--------", X"00010000", X"00020000"),

  ('1', "10010", "-----", "-----", X"00040000", X"--------", X"--------"),
  ('1', "10011", "-----", "-----", X"00080000", X"--------", X"--------"),
  ('0', "-----", "10010", "10011", X"--------", X"00040000", X"00080000"),

  ('1', "10100", "-----", "-----", X"00100000", X"--------", X"--------"),
  ('1', "10101", "-----", "-----", X"00200000", X"--------", X"--------"),
  ('0', "-----", "10100", "10101", X"--------", X"00100000", X"00200000"),

  ('1', "10110", "-----", "-----", X"00400000", X"--------", X"--------"),
  ('1', "10111", "-----", "-----", X"00800000", X"--------", X"--------"),
  ('0', "-----", "10110", "10111", X"--------", X"00400000", X"00800000"),

  ('1', "11000", "-----", "-----", X"01000000", X"--------", X"--------"),
  ('1', "11001", "-----", "-----", X"02000000", X"--------", X"--------"),
  ('0', "-----", "11000", "11001", X"--------", X"01000000", X"02000000"),

  ('1', "11010", "-----", "-----", X"04000000", X"--------", X"--------"),
  ('1', "11011", "-----", "-----", X"08000000", X"--------", X"--------"),
  ('0', "-----", "11010", "11011", X"--------", X"04000000", X"08000000"),

  ('1', "11100", "-----", "-----", X"10000000", X"--------", X"--------"),
  ('1', "11101", "-----", "-----", X"20000000", X"--------", X"--------"),
  ('0', "-----", "11100", "11101", X"--------", X"10000000", X"20000000"),

  ('1', "11110", "-----", "-----", X"40000000", X"--------", X"--------"),
  ('1', "11111", "-----", "-----", X"80000000", X"--------", X"--------"),
  ('0', "-----", "11110", "11111", X"--------", X"40000000", X"80000000")
  );

BEGIN

  UUT : ENTITY work.register_file GENERIC MAP (
    N => N,
    SIZE => SIZE
    )
    PORT MAP(
      clk => clk,
      wr_ena => sig.wr_ena,
      wr_sel => sig.wr_sel,
      rd_sel_1 => sig.rd_sel_1,
      rd_sel_2 => sig.rd_sel_2,
      wr => sig.wr,
      rd_1 => sig.rd_1,
      rd_2 => sig.rd_2
    );

  tick : PROCESS
  BEGIN
    clk <= '0';
    WAIT FOR TIME_SPAN / 2;
    clk <= '1';
    WAIT FOR TIME_SPAN / 2;
  END PROCESS;

  main : PROCESS
  BEGIN
    test_runner_setup(runner, runner_cfg);

    FOR i IN tests'RANGE LOOP

      sig.wr_ena <= tests(i).wr_ena;
      sig.wr_sel <= tests(i).wr_sel;
      sig.rd_sel_1 <= tests(i).rd_sel_1;
      sig.rd_sel_2 <= tests(i).rd_sel_2;
      sig.wr <= tests(i).wr;

      WAIT FOR TIME_SPAN;

      ASSERT (sig.rd_1 = tests(i).rd_1 OR tests(i).rd_1 = X"--------")
      REPORT "test " & INTEGER'image(i) & " failed [rd_1]" SEVERITY error;

      ASSERT (sig.rd_2 = tests(i).rd_2 OR tests(i).rd_2 = X"--------")
      REPORT "test " & INTEGER'image(i) & " failed [rd_2]" SEVERITY error;

    END LOOP;

    WAIT FOR TIME_SPAN;
    test_runner_cleanup(runner);
    WAIT;

  END PROCESS;

END tb;